module ALU_slt
(
  output result,
  input operandA,
  input operandB
);

endmodule
