`define AND and #330

module ALU_slt
(
  output result,
  input operandA,
  input operandB
);

endmodule
